`define REG_MY 0
`define REG_R1 1
`define REG_R2 2
`define REG_R3 3
`define REG_R4 4
`define REG_R5 5
`define REG_R6 6
`define REG_R7 7
`define REG_R8 8
`define REG_ZERO 9
`define REG_VIDEO 9
`define REG_X 10
`define REG_Y 11
`define REG_XMINUS 12
`define REG_XPLUS 13
`define REG_YMINUS 14
`define REG_YPLUS 15

`define LI 4'd0
`define UNL 4'd1
`define ADD 4'd2
`define SUB 4'd3
`define AND 4'd4
`define OR 4'd5
`define NOR 4'd6
`define SEQ 4'd7
`define SLT 4'd8
`define MUL 4'd9
`define SHR 4'd10
`define FMUL 4'd11
`define JUMP 4'd12
`define CALL 4'd13
`define RET 4'd14
